
typedef enum logic[3:0]{
    S0,  S1,  S2,  S3,  S4,
    S5,  S6,  S7,  S8,  S9,
    S10, S11, S12
} state_t;


parameter DELAY = 1;
parameter TRUE  = 1'b1;
parameter FALSE = 1'b0;